
module alu( in1 , in2 , opcode , out , flag );


endmodule
